** sch_path: /home/Joerdson/IHP-Open-PDK/ihp-sg13g2/libs.tech/xschem/LC_VCO.sch
**.subckt LC_VCO LO- LO+ VCC ICC GND VCTR
*.iopin LO-
*.iopin LO+
*.iopin VCC
*.iopin ICC
*.iopin GND
*.iopin VCTR
XMN3 LO+ LO- net1 GND sg13_lv_nmos w=40.0u l=0.13u ng=5 m=1
XMN4 LO- LO+ net1 GND sg13_lv_nmos w=40.0u l=0.13u ng=5 m=1
XMN1 ICC ICC GND GND sg13_lv_nmos w=120.0u l=0.13u ng=15 m=1
XMN12 net1 ICC GND GND sg13_lv_nmos w=120.0u l=0.13u ng=15 m=1
XC1 VCC LO+ cap_cmim w=8.73e-6 l=9.42e-6 m=1
XRp1 LO+ VCC rppd w=10.77e-6 l=8.92e-6 m=1 b=0
XC2 VCC LO- cap_cmim w=8.73e-6 l=9.42e-6 m=1
XRp2 LO- VCC rppd w=10.77e-6 l=8.92e-6 m=1 b=0
L1 VCC LO+ 2.006n m=1
L2 VCC LO- 2.006n m=1
XCvar LO+ VCTR LO- net1 sg13_hv_svaricap W=9.74e-6 L=0.8e-6 Nx=2
**.ends
.end
